module cordic
(
input clk,
input rst_n,
input [63:0] operand_1,
input [63:0] X_res, Y_res, Z_res,
input [3:0] state,
output reg [5:0] cordic_cnt,
output reg [63:0] Z_1, Z_2,       // the output to the add module
output reg [63:0] X_1, X_2, 
output reg [63:0] Y_1, Y_2
);

wire [63:0] atan_table [0:30];
wire [63:0] h_table [0:24];
reg [63:0] new_X_1, new_X_2;
reg [63:0] new_Y_1, new_Y_2;
reg [63:0] new_Z_1, new_Z_2;
reg [63:0] X_tmp, new_X_tmp;
reg [63:0] Y_tmp, new_Y_tmp;
reg [63:0] Z_tmp, new_Z_tmp;
reg need_repeated;
reg need_bias;

parameter IDLE = 4'd0, COMP = 4'd1, ADD = 4'd2, MUL = 4'd3, DIV = 4'd4, SIN_COS = 4'd5, SQUARE_ROOT = 4'd6, CORRECT_MODE = 4'd7, NATURAL_LOG = 4'd8;
integer i;

always @(posedge clk) begin
    if (~rst_n) begin
        cordic_cnt <= 0;
        X_1 <= 0;
        X_2 <= 0;
        Y_1 <= 0;
        Y_2 <= 0;
        Z_1 <= 0;
        Z_2 <= 0;
        need_repeated <= 0;
        X_tmp <= 0;
        Y_tmp <= 0;
        Z_tmp <= 0;
        need_bias <= 0;
    end
    else begin
        if (state == SIN_COS) begin
            if (cordic_cnt == 30)
                cordic_cnt <= 0;
            else
                cordic_cnt <= cordic_cnt + 1;
            X_1 <= new_X_1;
            X_2 <= new_X_2;
            Y_1 <= new_Y_1;
            Y_2 <= new_Y_2;
            Z_1 <= new_Z_1;
            Z_2 <= new_Z_2;
        end
        else if (state == SQUARE_ROOT) begin
            //need_bias <= new_need_bias;
            if (cordic_cnt == 30) begin
                cordic_cnt <= 0;
                need_repeated <= 0;
            end
            else if ((cordic_cnt == 4 || cordic_cnt == 13 || cordic_cnt == 40) && need_repeated == 0) begin
                cordic_cnt <= cordic_cnt;
                need_repeated <= 1;
            end
            else begin
                cordic_cnt <= cordic_cnt + 1;
                need_repeated <= 0;
            end

            X_1 <= new_X_1;
            X_2 <= new_X_2;
            Y_1 <= new_Y_1;
            Y_2 <= new_Y_2;
        end
        else if (state == NATURAL_LOG) begin
            if (cordic_cnt == 24) begin
                cordic_cnt <= 0;
                need_repeated <= 0;
                need_bias <= 0;
            end
            else if (cordic_cnt == 0 && need_bias == 0) begin
                cordic_cnt <= 0;
                need_bias <= 1;
            end
            else if (cordic_cnt <= 5 && need_repeated == 0 && need_bias == 1) begin
                cordic_cnt <= cordic_cnt;
                need_repeated <= 1;
            end
            else begin
                cordic_cnt <= cordic_cnt + 1;
                need_repeated <= 0;
            end
            X_1 <= new_X_1;
            X_2 <= new_X_2;
            X_tmp <= new_X_tmp;
            Y_1 <= new_Y_1;
            Y_2 <= new_Y_2;
            Y_tmp <= new_Y_tmp;
            Z_1 <= new_Z_1;
            Z_2 <= new_Z_2;
            Z_tmp <= new_Z_tmp;

        end
    end
end

always @* begin
    new_X_1 = 0;
    new_X_2 = 0;
    new_Y_1 = 0;
    new_Y_2 = 0;
    new_Z_1 = 0;
    new_Z_2 = 0;
    new_X_tmp = 0;
    new_Y_tmp = 0;
    new_Z_tmp = 0;

    if (state == SIN_COS) begin
        if (cordic_cnt == 0) begin
            new_X_1 = 64'b0011111111100011011011101001110111010111111011001011101110000000;   //0.607253
            new_X_2 = 0;

            new_Y_1 = 64'b0011111111100011011011101001110111010111111011001011101110000000;
            new_Y_2 = 0;

            new_Z_1 = operand_1;
            new_Z_2[63] = 1;
            new_Z_2[62:0] = atan_table[cordic_cnt][62:0];
        end
        else if (Z_res[63] == 0 || Z_res[62:0] == 0) begin
            new_X_1 = X_res;
            new_Y_1 = Y_res;
            new_Z_1 = Z_res;
            
            new_X_2[63] = ~Y_res[63];
            new_X_2[62:52] = Y_res[62:52] - cordic_cnt;
            new_X_2[51:0] = Y_res[51:0];

            new_Y_2[63:52] = X_res[63:52] - cordic_cnt;
            new_Y_2[51:0] = X_res[51:0];

            new_Z_2[63] = 1;
            new_Z_2[62:0]= atan_table[cordic_cnt][62:0];
        end
        else begin
            new_X_1 = X_res;
            new_Y_1 = Y_res;
            new_Z_1 = Z_res;

            new_X_2[63:52] = Y_res[63:52] - cordic_cnt;
            new_X_2[51:0] = Y_res[51:0];

            new_Y_2[63] = ~X_res[63];
            new_Y_2[62:52] = X_res[62:52] - cordic_cnt;
            new_Y_2[51:0] = X_res[51:0];

            new_Z_2 = atan_table[cordic_cnt];
        end
    end
    else if (state == SQUARE_ROOT) begin
        if (cordic_cnt == 0) begin
            new_X_1 = operand_1;
            new_X_2 = 64'b0011111111010000000000000000000000000000000000000000000000000000;

            new_Y_1 = operand_1;
            new_Y_2 = 64'b1011111111010000000000000000000000000000000000000000000000000000;
        end
        else begin
            if (Y_res[63] == 1) begin    // y < 0, di = 1
                new_X_1 = X_res;
                new_X_2[63] = Y_res[63];
                new_X_2[62:52] = Y_res[62:52] - cordic_cnt;
                new_X_2[51:0] = Y_res[51:0];

                new_Y_1 = Y_res;
                new_Y_2[63] = X_res[63];
                new_Y_2[62:52] = X_res[62:52] - cordic_cnt;
                new_Y_2[51:0] = X_res[51:0];
            end
            else begin
                new_X_1 = X_res;
                new_X_2[63] = ~Y_res[63];
                new_X_2[62:52] = Y_res[62:52] - cordic_cnt;
                new_X_2[51:0] = Y_res[51:0];

                new_Y_1 = Y_res;
                new_Y_2[63] = ~X_res[63];
                new_Y_2[62:52] = X_res[62:52] - cordic_cnt;
                new_Y_2[51:0] = X_res[51:0];
            end
        end
    end
    else if (state == NATURAL_LOG) begin
        if (cordic_cnt == 0 && need_bias == 0) begin
            new_X_1 = operand_1;
            new_X_2 = 64'b0011111111110000000000000000000000000000000000000000000000000000;

            new_Y_1 = operand_1;
            new_Y_2 = 64'b1011111111110000000000000000000000000000000000000000000000000000;

            new_Z_1 = 0;
            new_Z_2 = 0;
        end
        else if (cordic_cnt <= 5 && need_repeated == 0) begin   // retain value of Xres & Yres;
            new_X_tmp = X_res;
            new_Y_tmp = Y_res;
            new_Z_tmp = Z_res;

            new_X_1 = X_res;
            new_X_2[63] = ~X_res[63];
            new_X_2[62:52] = X_res[62:52] - (2 - cordic_cnt + 5);
            new_X_2[51:0] = X_res[51:0];

            new_Y_1 = Y_res;
            new_Y_2[63] = ~Y_res[63];
            new_Y_2[62:52] = Y_res[62:52] - (2 - cordic_cnt + 5);
            new_Y_2[51:0] = Y_res[51:0];

            new_Z_1 = 0;
            //new_Z_2 = h_table[cordic_cnt];
            new_Z_2 = 0;
        end
        else if (cordic_cnt <= 5 && need_repeated == 1) begin       
            if (X_tmp[63] == Y_tmp[63]) begin
                new_X_1 = X_tmp;
                new_X_2[63] = ~Y_res[63];
                new_X_2[62:0] = Y_res[62:0];

                new_Y_1 = Y_tmp;
                new_Y_2[63] = ~X_res[63];
                new_Y_2[62:0] = X_res[62:0];

                new_Z_1 = Z_tmp;
                new_Z_2 = h_table[cordic_cnt];
            end
            else begin
                new_X_1 = X_tmp;
                new_X_2 = Y_res;

                new_Y_1 = Y_tmp;
                new_Y_2 = X_res;

                new_Z_1 = Z_tmp;
                new_Z_2[63] = 1;
                new_Z_2[62:0] = h_table[cordic_cnt][62:0];
            end
        end
        else begin
            if (X_res[63] == Y_res[63]) begin
                new_X_1 = X_res;
                new_X_2[63] = ~Y_res[63];
                new_X_2[62:52] = Y_res[62:52] - (cordic_cnt - 5);
                new_X_2[51:0] = Y_res[51:0];

                new_Y_1 = Y_res;
                new_Y_2[63] = ~X_res[63];
                new_Y_2[62:52] = X_res[62:52] - (cordic_cnt - 5);
                new_Y_2[51:0] = X_res[51:0];

                new_Z_1 = Z_res;
                new_Z_2 = h_table[cordic_cnt];
            end
            else begin
                new_X_1 = X_res;
                new_X_2[63] = Y_res[63];
                new_X_2[62:52] = Y_res[62:52] - (cordic_cnt - 5);
                new_X_2[51:0] = Y_res[51:0];

                new_Y_1 = Y_res;
                new_Y_2[63] = X_res[63];
                new_Y_2[62:52] = X_res[62:52] - (cordic_cnt - 5);
                new_Y_2[51:0] = X_res[51:0];

                new_Z_1 = Z_res;
                new_Z_2[63] = 1;
                new_Z_2[62:0] = h_table[cordic_cnt][62:0];
            end
        end
    end
end

assign atan_table[0] = 64'b0100000001000110100000000000000000000000000000000000000000000000;  // 45       +5
assign atan_table[1] = 64'b0100000000111010100100001010011100110001101001100001110111000011;  // 26.5651
assign atan_table[2] = 64'b0100000000101100000100101000111010000000111110101110000000101110;  // 14.6262
assign atan_table[3] = 64'b0100000000011100100000000000010001001001001001111111111010000100;
assign atan_table[4] = 64'b0100000000001100100111000101010100110010011000010110010011010001;
assign atan_table[5] = 64'b0011111111111100101000110111100101001110010100101110001010100110;
assign atan_table[6] = 64'b0011111111101100101001010100001101010110001100110000111010110010;
assign atan_table[7] = 64'b0011111111011100101001011011010111101000010001001001111101110000;
assign atan_table[8] = 64'b0011111111001100101001011101001010001101110010101100100101000000;
assign atan_table[9] = 64'b0011111110111100101001011101100110110111001111000111000011001110;
assign atan_table[10] = 64'b0011111110101100101001011101101110000001100110011101110010101011;
assign atan_table[11] = 64'b0011111110011100101001011101101111110100001100010100011111100011;
assign atan_table[12] = 64'b0011111110001100101001011101110000010000110101110010001101000010;
assign atan_table[13] = 64'b0011111101111100101001011101110000011000000000001001101010101001;
assign atan_table[14] = 64'b0011111101101100101001011101110000011001110010101111011111110011;
assign atan_table[15] = 64'b0011111101011100101001011101110000011010001111011000011101100100;
assign atan_table[16] = 64'b0011111101001100101001011101110000011010010110100011010101011001;
assign atan_table[17] = 64'b0011111100111100101001011101110000011010011000010101111011010001;
assign atan_table[18] = 64'b0011111100101100101001011101110000011010011000110010100100101100;
assign atan_table[19] = 64'b0011111100011100101001011101110000011010011000111001101111000110;
assign atan_table[20] = 64'b0011111100001100101001011101110000011010011000111011100001101011;
assign atan_table[21] = 64'b0011111011111100101001011101110000011010011000111011111110010100;       // -16
assign atan_table[22] = 64'b0011111011101100101001011101110000011010011000111100000101011101;       // -17  
assign atan_table[23] = 64'b0011111011011100101001011101110000011010011000111100000111010001;
assign atan_table[24] = 64'b0011111011001100101001011101110000011010011000111100000111101101;
assign atan_table[25] = 64'b0011111010111100101001011101110000011010011000111100000111110100;
assign atan_table[26] = 64'b0011111010101100101001011101110000011010011000111100000111110111;
assign atan_table[27] = 64'b0011111010011100101001011101110000011010011000111100000111110111;
assign atan_table[28] = 64'b0011111010001100101001011101110000011010011000111100000111111001;
assign atan_table[29] = 64'b0011111001111100101001011101110000011010011000111100000111110101;
assign atan_table[30] = 64'b0011111001101100101001011101110000011010011000111100000111111000;
/*
assign atan_table[31] = 64'b0011111001011100101001011101110000011010011000111100000111111000; 
assign atan_table[32] = 64'b0011111001001100101001011101110000011010011000111100000111110101;  
assign atan_table[33] = 64'b0011111000111100101001011101110000011010011000111100000111111000;
assign atan_table[34] = 64'b0011111000101100101001011101110000011010011000111100000111111001;
assign atan_table[35] = 64'b0011111000011100101001011101110000011010011000111100000111110111;
assign atan_table[36] = 64'b0011111000001100101001011101110000011010011000111100000111111000;
assign atan_table[37] = 64'b0011110111111100101001011101110000011010011000111100000111111001;
assign atan_table[38] = 64'b0011110111101100101001011101110000011010011000111100000111110111;
assign atan_table[39] = 64'b0011110111011100101001011101110000011010011000111100000111110111;
assign atan_table[40] = 64'b0011110111001100101001011101110000011010011000111100000111111000;
assign atan_table[41] = 64'b0011110110111100101001011101110000011010011000111100000111111000;
assign atan_table[42] = 64'b0011110110101100101001011101110000011010011000111100000111110101;
assign atan_table[43] = 64'b0011110110011100101001011101110000011010011000111100000111111000;
assign atan_table[44] = 64'b0011110110001100101001011101110000011010011000111100000111111000;
assign atan_table[45] = 64'b0011110101111100101001011101110000011010011000111100000111111010;
assign atan_table[46] = 64'b0011110101101100101001011101110000011010011000111100000111111000;
assign atan_table[47] = 64'b0011110101011100101001011101110000011010011000111100000111110111;
assign atan_table[48] = 64'b0011110101001100101001011101110000011010011000111100000111111001;
assign atan_table[49] = 64'b0011110100111100101001011101110000011010011000111100000111110101;
assign atan_table[50] = 64'b0011110100101100101001011101110000011010011000111100000111111000;
assign atan_table[51] = 64'b0011110100011100101001011101110000011010011000111100000111110111;   
assign atan_table[52] = 64'b0011110100001100101001011101110000011010011000111100000111111010;        
assign atan_table[53] = 64'b0011110011111100101001011101110000011010011000111100000111111001;
assign atan_table[54] = 64'b0011110011101100101001011101110000011010011000111100000111111001;
assign atan_table[55] = 64'b0011110011011100101001011101110000011010011000111100000111110110;
assign atan_table[56] = 64'b0011110011001100101001011101110000011010011000111100000111111000;
assign atan_table[57] = 64'b0011110010111100101001011101110000011010011000111100000111111000;
assign atan_table[58] = 64'b00110100011001010010111011100001;
assign atan_table[59] = 64'b00110011111001010010111011100001;
assign atan_table[60] = 64'b00110011011001010010111011100001;
*/

assign h_table[0] = 64'b0100000000000110001010100100000011111101101000111110001111001100;   // idx = -5
assign h_table[1] = 64'b0100000000000011011000000111001010010100011000000010111001000011;
assign h_table[2] = 64'b0100000000000000100100101001000111101000111000110001100000011010;
assign h_table[3] = 64'b0011111111111011011110001100111001001000100100010010101101011001;
assign h_table[4] = 64'b0011111111110101101010100001011000111001010011010100100000011111;
assign h_table[5] = 64'b0011111111101111001000100111001010101110001100100101101001011010;  // idx = 0
assign h_table[6] = 64'b0011111111100001100100111110101001111010101011010000001100001100;  // idx = 1
assign h_table[7] = 64'b0011111111010000010110001010111011111010100000010001010001001011;
assign h_table[8] = 64'b0011111111000000000101011000100100011100100111101010111011110110;
assign h_table[9] = 64'b0011111110110000000001010101100010001010110100110111010110101100;
assign h_table[10] = 64'b0011111110100000000000010101010110001000100100011010111011100011;
assign h_table[11] = 64'b0011111110010000000000000101010101011000100010001010110011100000;
assign h_table[12] = 64'b0011111110000000000000000001010101010101100010001000100000101000;
assign h_table[13] = 64'b0011111101110000000000000000010101010101010110001000100101010011;
assign h_table[14] = 64'b0011111101100000000000000000000101010101010101011000110010010110;
assign h_table[15] = 64'b0011111101010000000000000000000001010101010101010101100010001001;
assign h_table[16] = 64'b0011111101000000000000000000000000010101010101010101010110001000;
assign h_table[17] = 64'b0011111100110000000000000000000000000101010101010101010101011001;
assign h_table[18] = 64'b0011111100100000000000000000000000000001010101010101010101010101;
assign h_table[19] = 64'b0011111100010000000000000000000000000000010101010101010101010101;
assign h_table[20] = 64'b0011111100000000000000000000000000000000000101010101010101010101;
assign h_table[21] = 64'b0011111011110000000000000000000000000000000001010101010101010110;
assign h_table[22] = 64'b0011111011100000000000000000000000000000000000010101010101010101;
assign h_table[23] = 64'b0011111011010000000000000000000000000000000000000101010101010100;
assign h_table[24] = 64'b0011111011000000000000000000000000000000000000000001010101010101;
/*
assign h_table[25] = 64'b0011111010110000000000000000000000000000000000000000010101010101;
assign h_table[26] = 64'b0011111010100000000000000000000000000000000000000000000101010101;
assign h_table[27] = 64'b0011111010010000000000000000000000000000000000000000000001010101;
assign h_table[28] = 64'b0011111010000000000000000000000000000000000000000000000000010101;
assign h_table[29] = 64'b0011111001110000000000000000000000000000000000000000000000000101;
*/
endmodule

